LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY sixty_counter IS
PORT(clk :IN STD_LOGIC; reset:IN STD_LOGIC;
 countl,countm :OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END sixty_counter;

ARCHITECTURE ar OF sixty_counter IS
SIGNAL l,m :INTEGER:=0;
SIGNAL lu,mu:UNSIGNED(3 DOWNTO 0);
BEGIN
PROCESS(clk,reset)
BEGIN
IF(reset ='0') THEN   
l<=0;
m<=0;
ELSIF(reset ='1') THEN   
   --counter is working
IF(clk'EVENT AND clk = '1') THEN
IF(m=5 AND l=9) THEN 
m <=m;
l <=l;
ELSIF(l=9) THEN
l <=0;
m <= m+1;
ELSE
l <= l+1;
END IF;
END IF;
END IF;

END PROCESS;
mu <= to_unsigned(m,4);
lu <= to_unsigned(l,4);
countl <= std_logic_vector(lu);
countm <= std_logic_vector(mu);
END ar ;



